
// -------------------------------- //
//	By: Bryce Keen	
//	Created: 08/13/2023
// -------------------------------- //
//	Last Modified: 08/13/2023

//
//	BEAN_2.v
//		The BEAN-2 is a RV32I implementation 
//    microarchitecture of the BEAN-2 follows a 5 stage pipelined CPU
//    with flush and stall capabilities
//    

// module BEAN_2 (clk, reset);


//   datapath data_unit(
//     .clk(clk), 
//     .reset(reset),
//     .reg_WE(reg_WE),
//     .rs1_SEL(rs1_SEL), 
//     .rs2_SEL(rs2_SEL),
//     .pc_SEL(pc_SEL), 
//     .reg_SEL(reg_SEL),
//     .imm_SEL(imm_SEL),
//     .ALU_SEL(ALU_SEL),
//     .Instr(Instr),
//     .memDataRD(memDataRD),
//     .pc(pc),
//     .memDataWD(memDataWD), 
//     .memAdrs(memAdrs),

//     .stall_F(stall_F), 
//     .stall_D(stall_D), 
//     .stall_E(stall_E), 
//     .stall_M(stall_M), 
//     .stall_WB(stall_WB),
//     .flush_F(flush_F), 
//     .flush_D(flush_D), 
//     .flush_E(flush_E), 
//     .flush_M(flush_M), 
//     .flush_WB(flush_WB));




//   control_logic control_unit(
//     .clk(clk), 
//     .reset(reset),
//     .opcode(opcode), 
//     .funct7(funct7), 
//     .funct3(funct3), 
//     .jump(jump), 
//     .ALU_SEL(ALU_SEL), 
//     .dmem_SEL(dmem_SEL), 
//     .imm_SEL(imm_SEL), 
//     .reg_SEL(reg_SEL), 
//     .pc_SEL(pc_SEL), 
//     .dmem_WE(dmem_WE), 
//     .reg_WE(reg_WE), 
//     .rs1_SEL(rs1_SEL), 
//     .rs2_SEL(rs2_SEL),

//     .stall_E(stall_E), 
//     .stall_M(stall_M), 
//     .stall_WB(stall_WB),
//     .flush_E(flush_E), 
//     .flush_M(flush_M), 
//     .flush_WB(flush_WB));


// // Hazard Unit




// endmodule


